module Gen_12ROT(input [3:0] k, output wire [17:0] Rre,
                                output wire [17:0] Rim);
  assign Rre = (k==0)? 65536 :  // cos(0π/6) * 2^16
               (k==1)? 56756 :  // cos(1π/6) * 2^16
               (k==2)? 32768 :  // cos(2π/6) * 2^16
               (k==3)? 0 :      // cos(3π/6) * 2^16
               (k==4)? -32768 : // cos(4π/6) * 2^16
               (k==5)? -56756 : // cos(5π/6) * 2^16
               (k==6)? -65536 : // cos(6π/6) * 2^16
               (k==7)? -56756 : // cos(7π/6) * 2^16
               (k==8)? -32768 : // cos(8π/6) * 2^16
               (k==9)? 0 :      // cos(9π/6) * 2^16
               (k==10)? 32768 : // cos(10π/6) *2^16
               (k==11)? 56756 : // cos(11π/6) *2^16
                       0 ;
  assign Rim = (k==0)? 0 :      // sin(0π/6) *2^16
               (k==1)? 32768 :  // sin(1π/6) *2^16
               (k==2)? 56756 :  // sin(2π/6) *2^16
               (k==3)? 65536 :  // sin(3π/6) *2^16
               (k==4)? 56756 :  // sin(4π/6) *2^16
               (k==5)? 32768 :  // sin(5π/6) *2^16
               (k==6)? 0 :      // sin(6π/6) *2^16
               (k==7)? -32768 : // sin(7π/6) *2^16
               (k==8)? -56756 : // sin(8π/6) *2^16
               (k==9)? -65536 : // sin(9π/6) *2^16
               (k==10)?-56756 : // sin(10π/6)*2^16
               (k==11)?-32768 : // sin(11π/6)*2^16
                       0 ;
endmodule